library verilog;
use verilog.vl_types.all;
entity Problem2BDF_vlg_vec_tst is
end Problem2BDF_vlg_vec_tst;
