library verilog;
use verilog.vl_types.all;
entity ALU_unit_vlg_vec_tst is
end ALU_unit_vlg_vec_tst;
