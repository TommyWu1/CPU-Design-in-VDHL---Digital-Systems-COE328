library verilog;
use verilog.vl_types.all;
entity Problem1BDF_vlg_vec_tst is
end Problem1BDF_vlg_vec_tst;
