library verilog;
use verilog.vl_types.all;
entity Problem3BDF_vlg_vec_tst is
end Problem3BDF_vlg_vec_tst;
